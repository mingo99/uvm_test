interface my_if(input clk, input rstn);

    logic [7:0] data;
    logic       valid;

endinterface: my_if